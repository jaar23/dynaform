module enums

pub enum DataType {
	string
	integer
	float
	boolean
	date
	datetime
} 