module enums

pub enum FormItemKind {
	input
	file_input
	hidden_input
	textarea
	checkbox
	radio
	selection
	label
	date_picker
	datetime_picker
	switch
}