module service

pub fn create() {
	println('create new form template')
}