module enums

pub enum TemplateStatus {
	dev
	prod
	archive
}